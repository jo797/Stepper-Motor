module stepper_rom (input clock, input [7:0] address,
			output reg [7:0] q);
//check the size of the address ??

			
endmodule
